// ------------------------------------------------------------------
// 4-bit ripple down counter (structural)
// ------------------------------------------------------------------

`include "DFlipFlop.v"
module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule

// ------------------------------------------------------------------
// 4-bit ripple down counter (dataflow)
// ------------------------------------------------------------------

`include "DFlipFlop.v"
module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule

// ------------------------------------------------------------------
// 4-bit ripple down counter (behavioral)
// ------------------------------------------------------------------

module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule

// ------------------------------------------------------------------
// 4-bit synchronous down counter (structural)
// ------------------------------------------------------------------

`include "TFlipFlop.v"
module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule

// ------------------------------------------------------------------
// 4-bit synchronous down counter (dataflow)
// ------------------------------------------------------------------

`include "TFlipFlop.v"
module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule

// ------------------------------------------------------------------
// 4-bit synchronous down counter (behavioral)
// ------------------------------------------------------------------

module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule

// ------------------------------------------------------------------
// 4-bit Johnson down counter (structural)
// ------------------------------------------------------------------

`include "DFlipFlop.v"
module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule

// ------------------------------------------------------------------
// 4-bit Johnson down counter (dataflow)
// ------------------------------------------------------------------

`include "DFlipFlop.v"
module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule

// ------------------------------------------------------------------
// 4-bit Johnson down counter (behavioral)
// ------------------------------------------------------------------

module counter(clk,out,reset_n);
	input clk,reset_n;
	output [3:0] out;
	
	// Implement counter here.
	
endmodule